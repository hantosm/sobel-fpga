module top(
    
);


endmodule